###############################################################################
#TSMC Library/IP Product
#Filename: tpb018v_3lm.lef
#Technology: 018
#Product Type: I/O PAD
#Product Name: tpb018v
#Version: 180a
###############################################################################
# 
#STATEMENT OF USE
#
#This information contains confidential and proprietary information of TSMC.
#No part of this information may be reproduced, transmitted, transcribed,
#stored in a retrieval system, or translated into any human or computer
#language, in any form or by any means, electronic, mechanical, magnetic,
#optical, chemical, manual, or otherwise, without the prior written permission
#of TSMC. This information was prepared for informational purpose and is for
#use by TSMC's customers only. TSMC reserves the right to make changes in the
#information at any time and without notice.
# 
###############################################################################

MACRO PAD80L
    CLASS BLOCK ;
    FOREIGN PAD80L 0.000 -72.500  ;
    ORIGIN 0.000 72.500 ;
    SIZE 80.000 BY 72.500 ;
    SYMMETRY X Y R90 ;
    OBS
        LAYER METAL1 ;
        RECT  0.000 -72.500 80.000 0.000 ;
        LAYER METAL2 ;
        RECT  0.000 -72.500 80.000 0.000 ;
        LAYER METAL3 ;
        RECT  0.000 -72.500 80.000 0.000 ;
    END
END PAD80L

MACRO PAD80L_OBV
    CLASS BLOCK ;
    FOREIGN PAD80L_OBV 0.000 -74.580  ;
    ORIGIN 0.000 74.580 ;
    SIZE 80.000 BY 74.580 ;
    SYMMETRY X Y R90 ;
    OBS
        LAYER METAL1 ;
        RECT  0.000 -74.580 80.000 0.000 ;
        LAYER METAL2 ;
        RECT  0.000 -74.580 80.000 0.000 ;
        LAYER METAL3 ;
        RECT  0.000 -74.580 80.000 0.000 ;
    END
END PAD80L_OBV

MACRO PAD80L_TRL
    CLASS BLOCK ;
    FOREIGN PAD80L_TRL 0.000 -72.500  ;
    ORIGIN 0.000 72.500 ;
    SIZE 80.000 BY 72.500 ;
    SYMMETRY X Y R90 ;
    OBS
        LAYER METAL1 ;
        RECT  0.000 -72.500 80.000 0.000 ;
        LAYER METAL2 ;
        RECT  0.000 -72.500 80.000 0.000 ;
        LAYER METAL3 ;
        RECT  0.000 -72.500 80.000 0.000 ;
    END
END PAD80L_TRL

END LIBRARY
